module RS485 #(clk_frequency)
(
    input clk,
    input rx,
    output tx
);

endmodule
