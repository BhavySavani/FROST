module uart #(parameter baud_rate,clk_frequency)
(
    input rx,
    input clk,
    output tx
);

endmodule 