module i2c#(parameter addr, clk_frequency)
(
    inout sda;
    output scl;
    input clk;
);

endmodule