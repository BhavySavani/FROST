module spi#(parameter clk_frequency)
(
    input clk,
    input miso,
    output mosi,
    output sclk,
    output cs
);

endmodule